//------------------------------------------------------------------------------
//
//  *** *** ***
// *   *   *   *
// *   *    *     Quantenna
// *   *     *    Connectivity
// *   *      *   Solutions
// * * *   *   *
//  *** *** ***
//     *
//------------------------------------------------------------------------------
`ifndef PKG_QCS_FIR_SV
`define PKG_QCS_FIR_SV

package qcs_dyn_pre_gen_pkg;
    import   uvm_pkg::*;
    import   qcs_gpio_pkg::*;
    `include "uvm_macros.svh"
    //
    `include "qcs_dyn_pre_gen_globals.svh"
    `include "qcs_dyn_pre_gen_cfg.sv"
    `include "qcs_dyn_pre_gen_item.sv"
    `include "qcs_dyn_pre_gen_sqr.sv"
    `include "qcs_dyn_pre_gen_drv.sv"
    `include "qcs_dyn_pre_gen_mon.sv"
    `include "qcs_dyn_pre_gen_ag.sv"
    
endpackage

`endif
