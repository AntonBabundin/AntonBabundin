//------------------------------------------------------------------------------
//
//  *** *** ***
// *   *   *   *
// *   *    *     Quantenna
// *   *     *    Connectivity
// *   *      *   Solutions
// * * *   *   *
//  *** *** ***
//     *
//------------------------------------------------------------------------------

package qcs_dyn_pre_gen_pkg_out;
    import   uvm_pkg::*;
    `include "uvm_macros.svh"
    //
    `include "qcs_dyn_pre_gen_globals_out.svh"
    `include "qcs_dyn_pre_gen_cfg_out.sv"
    `include "qcs_dyn_pre_gen_item_out.sv"
    `include "qcs_dyn_pre_gen_mon_out.sv"
    `include "qcs_dyn_pre_gen_ag_out.sv"
    
endpackage

