//------------------------------------------------------------------------------
//
//  *** *** ***
// *   *   *   *
// *   *    *     Quantenna
// *   *     *    Connectivity
// *   *      *   Solutions
// * * *   *   *
//  *** *** ***
//     *
//------------------------------------------------------------------------------
import  qcs_rst_gen_pkg::*;
import  qcs_clk_gen_pkg::*;
import  qcs_fir_pkg::*;
import  qcs_gpio_pkg::*;
