//------------------------------------------------------------------------------
//
//  *** *** ***
// *   *   *   *
// *   *    *     Quantenna
// *   *     *    Connectivity
// *   *      *   Solutions
// * * *   *   *
//  *** *** ***
//     *
//------------------------------------------------------------------------------
//---- sequences
`include  "base_sq.sv"
`include  "start_sq.sv"
`include  "tb_checkin_sq.sv"
`include  "fir_rx_zero_tst_sq.sv"
`include  "fir_rx_max_tst_sq.sv"
`include  "fir_rx_chirp_tst_sq.sv"
`include  "fir_rx_overflow_tst_sq.sv"


//---- tests
`include  "base_tst.sv"
`include  "start_tst.sv"
`include  "tb_checkin_tst.sv"
`include  "fir_rx_zero_tst.sv"
`include  "fir_rx_max_tst.sv"
`include  "fir_rx_chirp_tst.sv"
`include  "fir_rx_overflow_tst.sv"
