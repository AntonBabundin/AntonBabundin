//------------------------------------------------------------------------------
//
//  *** *** ***
// *   *   *   *
// *   *    *     Quantenna
// *   *     *    Connectivity
// *   *      *   Solutions
// * * *   *   *
//  *** *** ***
//     *
//------------------------------------------------------------------------------
`ifndef PKG_QCS_CHKP_PROBE_SV
`define PKG_QCS_CHKP_PROBE_SV

package qcs_chkp_probe_pkg;
  import   uvm_pkg::*;
  `include "uvm_macros.svh"
  //----
  `include "qcs_chkp_probe_globals.svh"
endpackage

`endif
